module icache#(
  localparam ICACHE_NUM_ASSOCIATE = 4,
  localparam ICACHE_OFFSET_WIDTH  = 8,
  localparam ICACHE_INDEX_WIDTH   = 8,
  localparam ICACHE_TAG_WIDTH     = 8
)(
  input logic  clk_i,
  input logic  icache_req_i,
  output logic icache_ready_o,
  input logic  icache_req_vaddr_i,
  input logic  icache_req_paddr_i,
  output logic icache_resp_data_o
);






endmodule